library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ADT7420 is
    port (
        clk   : in std_logic;
        reset : in std_logic;
        
    );
end entity ADT7420;

architecture ADT7420_arch of ADT7420 is

begin

    

end architecture ADT7420_arch;
